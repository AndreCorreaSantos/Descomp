library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13; -- Instrucoes de 13 bits
          addrWidth: natural := 3 -- so preciso de 3 bits 
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0) -- 12 downto 0
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

    constant NOP  : std_logic_vector(3 downto 0) := "0000";
    constant LDA  : std_logic_vector(3 downto 0) := "0001";
    constant SOMA : std_logic_vector(3 downto 0) := "0010";
    constant SUB  : std_logic_vector(3 downto 0) := "0011";
    constant LDI : std_logic_vector(3 downto 0) := "0100";
    constant STA : std_logic_vector(3 downto 0) := "0101";
    
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
        tmp(0) := LDI & "000000100";
        tmp(1) := STA & "100000001";
        tmp(2) := LDI & "000000011";
        tmp(3) := STA & "100000000";
        tmp(4) := SOMA & "100000000";
        tmp(5) := SOMA & "100000000";
        tmp(6) := SOMA & "100000000";
        tmp(6) := SUB & "100000001";
        tmp(7) := NOP & "000000000";

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;